library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity alu is 
	port( X,Y : in std_logic_vector(15 downto 0);
		x0,x1 : in std_logic ;
		C_in: in std_logic;
		C_out, Z_out: out std_logic;
		S : out std_logic_vector(15 downto 0));
end entity;

architecture alu_behave of alu is
	signal sig1,sig2,sig3: std_logic_vector(15 downto 0);
	signal car1, car2 : std_logic;

	component SixteenBitAdder is
		port(x,y: in std_logic_vector(15 downto 0);
			z: out std_logic_vector(15 downto 0);
			car_in: in std_logic;
			car_out: out std_logic);
	end component;

	component SixteenBitSub is
		port(x,y: in std_logic_vector(15 downto 0);
			z: out std_logic_vector(15 downto 0);
			bor_in: in std_logic;
			bor_out: out std_logic);	
	end component;

	component SixteenBitNand is
		port(x,y: in std_logic_vector(15 downto 0);
			z: out std_logic_vector(15 downto 0));
	end component;

begin
	a: SixteenBitAdder port map (x => X, y => Y, z => sig1, car_in => C_in, car_out => car1);
	b: SixteenBitSub port map (x => X, y => Y, z => sig2, bor_in => C_in, bor_out => car2);
	c: SixteenBitNand port map (x => X, y => Y, z => sig3);

	process (x0, x1, sig1, sig2, sig3, car1, car2)
	begin
		if (x0 = '1' and x1 = '1') then
			S <= sig1; -- ADD operation
			C_out <= car1;
			Z_out <= not (sig1(0) and sig1(1) and sig1(2) and sig1(3) and sig1(4) and sig1(5) and sig1(6) and sig1(7) and sig1(8) and sig1(9) and sig1(10) and sig1(11) and sig1(12) and sig1(13) and sig1(14) and sig1(15));
		elsif (x0 = '1' and x1 = '0') then
			S <= sig2; -- SUB operation
			C_out <= car2;
			Z_out <= not (sig2(0) and sig2(1) and sig2(2) and sig2(3) and sig2(4) and sig2(5) and sig2(6) and sig2(7) and sig2(8) and sig2(9) and sig2(10) and sig2(11) and sig2(12) and sig2(13) and sig2(14) and sig2(15));
		elsif (x0 = '0' and x1 = '1') then
			S <= sig3; -- NAND operation
			C_out <= C_in;
			Z_out <= not (sig3(0) and sig3(1) and sig3(2) and sig3(3) and sig3(4) and sig3(5) and sig3(6) and sig3(7) and sig3(8) and sig3(9) and sig3(10) and sig3(11) and sig3(12) and sig3(13) and sig3(14) and sig3(15));
		end if;
	end process;

end alu_behave;